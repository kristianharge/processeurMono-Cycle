library IEEE;
use IEEE.STD_LOGIC_1164.all;
USE ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity EDS_TB is
 port( OK: out boolean:=FALSE);
end entity EDS_TB;

architecture BENCH of EDS_TB is
  constant TN: positive := 16;
  signal TA: std_logic_vector (TN-1 downto 0);
  signal TS: std_logic_vector(31 downto 0);
  
  component EDS is
    generic ( N: positive range 1 to 32);
    
    PORT(
		A :  IN  std_logic_vector (N-1 downto 0);
		S :  OUT  std_logic_vector (31 downto 0)
	);
  end component;
  
begin
  
  UUT: COMPONENT EDS
  generic map(
    N => TN
    )
    
  PORT MAP(
	  A => TA,
    S => TS
  );

  stimulus:process
  begin
        
        wait for 1 ns;
        TA <= "0000000000000001";
        wait for 1 ns;
        ASSERT signed(TS) /= signed(TA)REPORT "ERROR: EDS TEST 1 FAILED)" -- EDS Test 1
        SEVERITY FAILURE; 
        REPORT "EDS Test 1 passed." SEVERITY note;

        wait for 1 ns;
        TA <= "1111111111111001";
        wait for 1 ns;
        ASSERT signed(TS) /= signed(TA)REPORT "ERROR: EDS TEST 1 FAILED)" -- EDS Test 1
        SEVERITY FAILURE; 
        REPORT "EDS Test 1 passed." SEVERITY note;

        REPORT "Bench test is successfully finished." SEVERITY note;
        OK <= TRUE; -- La fin du banc de teste. Le r�sultat est bon.
        WAIT; -- Boucle infinie
  end process;

  
end architecture BENCH;

